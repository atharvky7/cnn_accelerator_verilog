// Parameter include file for CNN accelerator
